module empty ();
endmodule
module empty2 ;
endmodule

