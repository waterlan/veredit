module test (a, b, c, d, e, f);

  i1 buf (.z(d), .a(c));
assign a = b;
output d;
input [2:0] f;
output [2:0] e;
wire a;
  i0 buf (.z(d), .a(c));
assign e = f;
input c;

wire d;

output a;
input b ;

endmodule

