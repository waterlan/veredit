
module test1 ( Z, A,B );
output Z;
input  A;
input  B;

wire a ;
wire [1:0] b, bb;
wire [2:0] bbb;
wire c, d;
supply0  zero, zero2;
tri TT;


endmodule

module test2 ( Z, A,B );
output Z;
input  A;
input  B;

wire a ;
wire [1:0] b;
wire c, d;


endmodule

