module a (z, a);
input a;
output z;

assign z = a;

endmodule

module b (z, a);
input a;
output z;

assign z = a;

endmodule

module c (z, a);
input a;
output z;

assign z = a;

endmodule

module d (z, a);
input a;
output z;

assign z = a;

endmodule

